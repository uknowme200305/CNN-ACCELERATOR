module reg_block#(parameter WIDTH = 8)(input clk , rst , en , input [WIDTH -1:0]d , output reg [WIDTH -1:0]q);

always@(posedge clk or posedge rst)begin 
    if(rst)
        q<=0;
        else if(en)
        q<=d;
end

endmodule